`timescale 1ns / 1ps

module SSD(D,C ,B);
    parameter N=4;
    output [6:0] D;
    output [6:0] C;
    input [3:0] B;
    //reg [N-1:0] B;
    reg [6:0] C;
    reg [6:0] D;
always @(B,C)
    begin
    case (B)
        4'b0000: C=7'b1000000;
        4'b0001: C=7'b1111001;
        4'b0010: C=7'b0100100;
        4'b0011: C=7'b0110000;
        4'b0100: C=7'b0011001;
        4'b0101: C=7'b0010010;
        4'b0110: C=7'b0000010;
        4'b0111: C=7'b1111000;
        4'b1000: C=7'b0000000;
        4'b1001: C=7'b1111000;
        4'b1010: C=7'b0000010;
        4'b1011: C=7'b0010010;
        4'b1100: C=7'b0011001;
        4'b1101: C=7'b0110000;
        4'b1110: C=7'b0100100;
        4'b1111: C=7'b1111001;
        endcase
   case (B)
        4'b0000: D=7'b1111111;
        4'b0001: D=7'b1111111;
        4'b0010: D=7'b1111111;
        4'b0011: D=7'b1111111;
        4'b0100: D=7'b1111111;
        4'b0101: D=7'b1111111;
        4'b0110: D=7'b1111111;
        4'b0111: D=7'b1111111;
        4'b1000: D=7'b0111111;
        4'b1001: D=7'b0111111;
        4'b1010: D=7'b0111111;
        4'b1011: D=7'b0111111;
        4'b1100: D=7'b0111111;
        4'b1101: D=7'b0111111;
        4'b1110: D=7'b0111111;
        4'b1111: D=7'b0111111;
        endcase
  end 
endmodule
